`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:50:36 07/25/2021 
// Design Name: 
// Module Name:    partialproduct16bit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module partial16bit(x,y,a0,a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12,a13,a14,a15);
 input [15:0]x,y;
 output [15:0]a0,a1,a2,a3,a4,a5,a6,a7,a8,a9,a10;
 output [15:0]a11,a12,a13,a14,a15;
 
 assign a0= {x[0]&y[15],x[0]&y[14],x[0]&y[13],x[0]&y[12],x[0]&y[11],x[0]&y[10], x[0]&y[9],x[0]&y[8],x[0]&y[7],x[0]&y[6],x[0]&y[5],x[0]&y[4],x[0]&y[3],x[0]&y[2], x[0]&y[1],x[0]&y[0]};
 assign a1={x[1]&y[15],x[1]&y[14],x[1]&y[13],x[1]&y[12],x[1]&y[11],x[1]&y[10], x[1]&y[9],x[1]&y[8],x[1]&y[7],x[1]&y[6],x[1]&y[5],x[1]&y[4],x[1]&y[3],x[1]&y[2], x[1]&y[1],x[1]&y[0]};
 assign a2={x[2]&y[15],x[2]&y[14],x[2]&y[13],x[2]&y[12],x[2]&y[11],x[2]&y[10], x[2]&y[9],x[2]&y[8],x[2]&y[7],x[2]&y[6],x[2]&y[5],x[2]&y[4],x[2]&y[3],x[2]&y[2], x[2]&y[1],x[2]&y[0]};
 assign a3={x[3]&y[15],x[3]&y[14],x[3]&y[13],x[3]&y[12],x[3]&y[11],x[3]&y[10], x[3]&y[9],x[3]&y[8],x[3]&y[7],x[3]&y[6],x[3]&y[5],x[3]&y[4],x[3]&y[3],x[3]&y[2], x[3]&y[1],x[3]&y[0]};
 assign a4={x[4]&y[15],x[4]&y[14],x[4]&y[13],x[4]&y[12],x[4]&y[11],x[4]&y[10], x[4]&y[9],x[4]&y[8],x[4]&y[7],x[4]&y[6],x[4]&y[5],x[4]&y[4],x[4]&y[3],x[4]&y[2], x[4]&y[1],x[4]&y[0]};
 assign a5={x[5]&y[15],x[5]&y[14],x[5]&y[13],x[5]&y[12],x[5]&y[11],x[5]&y[10], x[5]&y[9],x[5]&y[8],x[5]&y[7],x[5]&y[6],x[5]&y[5],x[5]&y[4],x[5]&y[3],x[5]&y[2], x[5]&y[1],x[5]&y[0]};
 assign a6={x[6]&y[15],x[6]&y[14],x[6]&y[13],x[6]&y[12],x[6]&y[11],x[6]&y[10], x[6]&y[9],x[6]&y[8],x[6]&y[7],x[6]&y[6],x[6]&y[5],x[6]&y[4],x[6]&y[3],x[6]&y[2], x[6]&y[1],x[6]&y[0]};
 assign a7={x[7]&y[15],x[7]&y[14],x[7]&y[13],x[7]&y[12],x[7]&y[11],x[7]&y[10], x[7]&y[9],x[7]&y[8],x[7]&y[7],x[7]&y[6],x[7]&y[5],x[7]&y[4],x[7]&y[3],x[7]&y[2], x[7]&y[1],x[7]&y[0]};
 assign a8={x[8]&y[15],x[8]&y[14],x[8]&y[13],x[8]&y[12],x[8]&y[11],x[8]&y[10], x[8]&y[9],x[8]&y[8],x[8]&y[7],x[8]&y[6],x[8]&y[5],x[8]&y[4],x[8]&y[3],x[8]&y[2], x[8]&y[1],x[8]&y[0]};
 assign a9={x[9]&y[15],x[9]&y[14],x[9]&y[13],x[9]&y[12],x[9]&y[11],x[9]&y[10], x[9]&y[9],x[9]&y[8],x[9]&y[7],x[9]&y[6],x[9]&y[5],x[9]&y[4],x[9]&y[3],x[9]&y[2], x[9]&y[1],x[9]&y[0]};
 assign a10={x[10]&y[15],x[10]&y[14],x[10]&y[13],x[10]&y[12],x[10]&y[11],x[10]&y[10], x[10]&y[9],x[10]&y[8],x[10]&y[7],x[10]&y[6],x[10]&y[5],x[10]&y[4],x[10]&y[3],x[10]&y[2], x[10]&y[1],x[10]&y[0]};
 assign a11={x[11]&y[15],x[11]&y[14],x[11]&y[13],x[11]&y[12],x[11]&y[11],x[11]&y[10], x[11]&y[9],x[11]&y[8],x[11]&y[7],x[11]&y[6],x[11]&y[5],x[11]&y[4],x[11]&y[3],x[11]&y[2], x[11]&y[1],x[11]&y[0]};
assign a12={x[12]&y[15],x[12]&y[14],x[12]&y[13],x[12]&y[12],x[12]&y[11],x[12]&y[10], x[12]&y[9],x[12]&y[8],x[12]&y[7],x[12]&y[6],x[12]&y[5],x[12]&y[4],x[12]&y[3],x[12]&y[2], x[12]&y[1],x[12]&y[0]};
assign a13={x[13]&y[15],x[13]&y[14],x[13]&y[13],x[13]&y[12],x[13]&y[11],x[13]&y[10], x[13]&y[9],x[13]&y[8],x[13]&y[7],x[13]&y[6],x[13]&y[5],x[13]&y[4],x[13]&y[3],x[13]&y[2], x[13]&y[1],x[13]&y[0]};
assign a14={x[14]&y[15],x[14]&y[14],x[14]&y[13],x[14]&y[12],x[14]&y[11],x[14]&y[10], x[14]&y[9],x[14]&y[8],x[14]&y[7],x[14]&y[6],x[14]&y[5],x[14]&y[4],x[14]&y[3],x[14]&y[2], x[14]&y[1],x[14]&y[0]};
assign a15={x[15]&y[15],x[15]&y[14],x[15]&y[13],x[15]&y[12],x[15]&y[11],x[15]&y[10], x[15]&y[9],x[15]&y[8],x[15]&y[7],x[15]&y[6],x[15]&y[5],x[15]&y[4],x[15]&y[3],x[15]&y[2], x[15]&y[1],x[15]&y[0]};
  
  endmodule







